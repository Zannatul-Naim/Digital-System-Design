module nand_gate(y, a, b);
  
    input a, b;
    output y;
    nand(y, a, b);
  
endmodule
