module xor_gate(output y, input a, input b);  
    xnor(y, a, b);
  
endmodule
