module and_gate(y, a, b);
  
    input a, b;
    output y;
    and(y, a, b);
  
endmodule
