module not_gate(output y, input x);
  
  not(y, x);
  
endmodule
