module xor_gate(output y, input a, input b);
  
    xor(y, a, b);
  
endmodule
