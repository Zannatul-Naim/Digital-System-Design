module or_gate(y, a, b); 
    input a, b;
    output y;
    nor(y, a, b);  
  
endmodule
